module JAM (
    input CLK,
    input RST,
    output [3:0] MatchCount,
    output [9:0] MinCost,
    output       Valid,

    output [2:0] W,
    output [2:0] J,
    input  [6:0] Cost
);



endmodule


